module bit_a(input a, input b, output logic c)
    assign c = a + b;
endmodule