module hello;
  initial 
    $display("Hello World");
endmodule
